library ieee;
use ieee.std_logic_1164.all;

entity One_Bit_Adder is
  port ( a: in std_logic;
         b: in std_logic;
         c: in std_logic;
         d: out std_logic;
         e: out std_logic
       );
     end One_Bit_Adder;
     
  architecture struct of One_Bit_Adder is
  
    component AND_gate is
      port ( x: in std_logic;
             y: in std_logic;
             z: out std_logic
           );
      end component;
      
    component OR_gate is
      port ( x: in std_logic;
             y: in std_logic;
             z: out std_logic
           );
      end component;            
      
    component XOR_gate is
      port ( a: in std_logic;
             b: in std_logic;
             c: out std_logic
           );
      end component;
      
      signal temp1: std_logic;
      signal temp2: std_logic;
      signal temp3: std_logic;
      
      begin
        
        --map signals
        map_XOR_gate: XOR_gate port map (a, b, temp1);
        map_XOR_gate2: XOR_gate port map (temp1, c, d);
        map_AND_gate: AND_gate port map (a, b, temp2);
        map_AND_gate2: AND_gate port map (temp1, c, temp3);
        map_OR_gate: OR_gate port map (temp2, temp3, e);
          
        end struct;